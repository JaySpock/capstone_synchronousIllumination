library IEEE;
use IEEE.STD_LOGIC_1164.ALL; 
use IEEE.NUMERIC_STD.ALL; 
use IEEE.std_logic_unsigned.all; 

LIBRARY altera; 
USE altera.altera_primitives_components.all;
  

entity project is 

    port(   clk    			: in std_logic; 										-- Clock signal

            KEY    			: in std_logic;										-- Startup switch
				
				DATA 	 			: in std_logic;										-- Current bit from Camera
				
				DATA_OUT 		: out std_logic;										-- Rising edge indicates EOF
				
				LED_OUT			: out std_logic_vector(2 downto 0);				-- LED output for the pins--
				
            LED    			: out std_logic_vector(2 downto 0)); 			-- LED output for development board LEDs

end entity; 

  

architecture blink_arch of project is 

	component datacapture
	port(
		 clk: in std_logic;
		 clk_enable: in std_logic;
		 ready_to_capture: out std_logic;
		 Data_out: in std_logic_vector(4 downto 0); 
		 Calibration: in std_logic; 
		 New_Frame: in std_logic); 
	end component;


	signal FIFO_reg		: std_logic_vector(61 downto 0) := "11111111111111111111111111111111111111111111111111111111111111";

	signal LED_output 	: std_logic_vector(2 downto 0) := "110"; -- RED?
	
	signal LED_BUFFER 	: std_logic := '1'; 
	
	signal NEW_FRAME		: std_logic := '0'; 
	
	signal Calibration	: std_logic := '0'; 
	
	signal DATA_BUFFER	: std_logic;

	signal cnt         	: INTEGER RANGE 0 TO 25000000;

	signal startup_frame	: INTEGER RANGE 0 to 9 := 4;
	
	signal cal_cnt			: INTEGER RANGE 0 to 2;

	begin 
	
		u0: datacapture
			port map(clk=>clk,
						clk_enable=>'1',
						Data_out=>(Calibration & NEW_FRAME & LED_output),
						Calibration=>Calibration,
						New_Frame=>NEW_FRAME);
						
		DATA_OUT <= NEW_FRAME;

		LED<= LED_output; 
		
		LED_out <= LED_output;
		
--	process(KEY)
--		begin
--			if(KEY = '1') then
--				startup_frame <= 0;
--			end if;
--	end process;
--				
	 process (clk)
			begin
			
				if (rising_edge(clk)) then	
				
					if (DATA_BUFFER = '1') then
				
						cnt <= cnt + 1;
						
					end if;
					
					for address in 61 downto 1 loop
						
						FIFO_reg(address) <= FIFO_reg(address - 1);
							
					end loop;
				
--						
					FIFO_reg(0) <= DATA;
					
--					FIFO_reg <= FIFO_reg(126 downto 0) & DATA;
					
					if(KEY = '0') then
							startup_frame <= 0;
					end if;
--					
					if (FIFO_reg = "00000000000000000000000000000000000000000000000000000000000000" and DATA_BUFFER = '0') then
					
						LED_BUFFER    <= LED_output(2);
					
						NEW_FRAME <= '1';
						DATA_BUFFER <= '1';
						cnt <= 0;
						
						case startup_frame is
							when 0	=> 
								Calibration <= '1';
								LED_output <= "111";						--NO LIGHT startup frame
								if(cal_cnt = 2) then
									startup_frame <= 1;
									cal_cnt <= 0;
								else
									cal_cnt <= cal_cnt + 1;
								end if;
								
							when 1	=>
--								LED_output <= "110";						--RED startup frame
								if(cal_cnt = 1) then
									LED_output <= "111";
									cal_cnt <= cal_cnt + 1;	
								elsif(cal_cnt = 0) then
									LED_output <= "110";
									cal_cnt <= cal_cnt + 1;	
								else
									LED_output <= "111";	
									startup_frame <= 2;
									cal_cnt <= 0;	
								end if;
	
							when 2	=>
								if(cal_cnt = 1) then
									LED_output <= "111";
									cal_cnt <= cal_cnt + 1;	
								elsif(cal_cnt = 0) then
									LED_output <= "101";
									cal_cnt <= cal_cnt + 1;	
								else
									LED_output <= "111";	
									startup_frame <= 3;
									cal_cnt <= 0;	
								end if;
	
							
--								LED_output <= "011";						--GREEN startup frame?
--								if(cal_cnt = 2) then
--									startup_frame <= 3;
--									cal_cnt <= 0;
--								else
--									cal_cnt <= cal_cnt + 1;
--								end if;
								
							when 3 	=>
								if(cal_cnt = 1) then
									LED_output <= "111";
									cal_cnt <= cal_cnt + 1;	
								elsif(cal_cnt = 0) then
									LED_output <= "011";
									cal_cnt <= cal_cnt + 1;	
								else
									LED_output <= "111";	
									startup_frame <= 4;
									cal_cnt <= 0;	
								end if;
								
--								LED_output <= "101";						--BLUE startup frame?
--								if(cal_cnt = 2) then
--									startup_frame <= 4;
--									cal_cnt <= 0;
--								else
--									cal_cnt <= cal_cnt + 1;
--								end if;
--								
							when others =>
								Calibration <= '0';
								case LED_output is
									when "110" =>
										LED_output <= "101";
									when "101" =>
										LED_output <= "011";
									when "011" =>
										LED_output <= "110";	
									when "111" =>
										LED_output <= "110";	
									when others =>
										LED_output <= "111";
--								LED_BUFFER    <= LED_output(2);
--								LED_output(2) <= LED_output(1);
--								LED_output(1) <= LED_output(0);
--								LED_output(0) <= LED_BUFFER;
								end case;						
						end case;
					elsif (DATA_BUFFER = '1' and cnt >25000) then
					
						NEW_FRAME <= '0';
						DATA_BUFFER <= '0';
						cnt <= 0;
					end if;
				end if;
			end process;
	end architecture; 


--library IEEE; 
--
--use IEEE.STD_LOGIC_1164.ALL; 
--
--use IEEE.NUMERIC_STD.ALL; 
--
--use IEEE.std_logic_unsigned.all; 
--
--  
--
--LIBRARY altera; 
--
--USE altera.altera_primitives_components.all; 
--
--  
--
--  
--
--entity project is 
--
--    port(    clk    : in std_logic; 
--
--            KEY    : in std_logic; 
--				
----				Vout	 : out std_logic;
--				
--				DATA 	 : in std_logic;
--				
--				DATA_OUT : out std_logic;
--				
--				LED_DATA_OUT : out std_logic_vector(2 downto 0);
--				
--            LED    : out std_logic_vector(2 downto 0)); 
--
--end entity; 
--
--  
--
--architecture blink_arch of project is 
--
--  
--
--	signal LED_output : std_logic_vector(2 downto 0) := "110"; 
--	
--	signal LED_BUFFER : std_logic; 
--	
--	signal word  :	std_logic_vector(11 downto 0);
--	
--	signal DATA_BUFFER : std_logic;
--
--	signal cnt         : INTEGER RANGE 0 TO 25000000;
--
--	type RW_type is array (0 to 15) of std_logic;
--
--	signal RW : RW_type;
--	
--  
--
--	begin 
--
--		
--
--		LED<= LED_output; 
--
--		LED_DATA_OUT <= LED_output;
--		
--		
--		
--	 process (clk)
--			begin
--			
--				if (clk'event and clk='1') then	
--				
--			
--					cnt <= cnt + 1;
--							
----					LED_output(3 downto 0) <= not LED_output(3 downto 0);
----					DATA_OUT <= DATA;
--					
--					for address in 15 downto 1 loop
--						
--						RW(address) <= RW(address - 1);
--							
--					end loop;
--				
----						
--					RW(0) <= DATA;
--					
--					word <= (RW(0) & RW(1) & RW(2) & RW(3) & RW(4) & RW(5) & RW(6) & RW(7) & RW(8) & RW(9) & RW(10) & RW(11));
--					
--					if (word = "000000000000" and DATA_BUFFER ='0') then
--					
--						DATA_OUT <= '1';
--						LED_BUFFER <= LED_output(2);
--						LED_output(2) <= LED_output(1);
--						LED_output(1) <= LED_output(0);
--						LED_output(0) <= LED_BUFFER;
--						DATA_BUFFER <= '1';
--						cnt <= 0;
--					
--					elsif (DATA_BUFFER = '1' and cnt >25000) then
--					
--						DATA_OUT <= '0';
--						DATA_BUFFER <= '0';
--						cnt <= 0;
--					end if;
--					
--				end if;
--			end process;
--
--
	  

--	end architecture; 
	component nios_setup is
		port (
			clk_clk                           : in  std_logic                    := 'X';             -- clk
			led_external_connection_export    : in  std_logic_vector(4 downto 0) := (others => 'X'); -- export
			reset_reset_n                     : in  std_logic                    := 'X';             -- reset_n
			switch_external_connection_export : out std_logic_vector(2 downto 0)                     -- export
		);
	end component nios_setup;

	u0 : component nios_setup
		port map (
			clk_clk                           => CONNECTED_TO_clk_clk,                           --                        clk.clk
			led_external_connection_export    => CONNECTED_TO_led_external_connection_export,    --    led_external_connection.export
			reset_reset_n                     => CONNECTED_TO_reset_reset_n,                     --                      reset.reset_n
			switch_external_connection_export => CONNECTED_TO_switch_external_connection_export  -- switch_external_connection.export
		);

